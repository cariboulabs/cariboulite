module complex_fifo #(
    parameter ADDR_WIDTH = 8,
    parameter DATA_WIDTH = 16
)
(
    input wire 			            wr_rst_i,
    input wire 			            wr_clk_i,
    input wire 			            wr_en_i,
    input wire [2*DATA_WIDTH-1:0]	wr_data_i,

    input wire 			            rd_rst_i,
    input wire 			            rd_clk_i,
    input wire 			            rd_en_i,
    output reg [2*DATA_WIDTH-1:0]	rd_data_o,

    output reg 			full_o,
    output reg 			empty_o
);

reg [ADDR_WIDTH-1:0]	wr_addr;
reg [ADDR_WIDTH-1:0]	rd_addr;

always @(posedge wr_clk_i) begin
    if (wr_rst_i) begin
        wr_addr <= 0;
        full_o <= 1'b0;
    end else begin
        if (wr_en_i) begin
            wr_addr <= wr_addr + 1'b1;
            full_o <= (wr_addr + 2) == rd_addr;
            mem_i[wr_addr] <= wr_data_i[31:16];
            mem_q[wr_addr] <= wr_data_i[15:0];
        end else begin
            full_o <= full_o & ((wr_addr + 1'b1) == rd_addr);
        end
    end
end

always @(posedge rd_clk_i) begin
    if (rd_rst_i) begin
        rd_addr <= 0;
        empty_o <= 1'b1;
    end else begin
        if (rd_en_i) begin
            rd_addr <= rd_addr + 1'b1;
            empty_o <= (rd_addr + 1) == wr_addr;
            rd_data_o[31:16] <= mem_i[rd_addr];
            rd_data_o[15:0] <= mem_q[rd_addr];
        end else begin
            empty_o <= empty_o & (rd_addr == wr_addr);
        end
    end
end

reg [DATA_WIDTH-1:0] mem_i[(1<<ADDR_WIDTH)-1:0];
reg [DATA_WIDTH-1:0] mem_q[(1<<ADDR_WIDTH)-1:0];

endmodule

// generate dual clocked memory
/*SB_RAM40_4K #(
    .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .WRITE_MODE(0),
    .READ_MODE(0)
) ram256x16_i_inst (
    .RDATA(rd_data_o[31:16]),
    .RADDR(rd_addr),
    .RCLK(rd_clk_i),
    .RCLKE(1),    //<<
    .RE(rd_en_i),
    .WADDR(wr_addr),
    .WCLK (wr_clk_i),
    .WCLKE(wr_en_i),    //<<
    .WDATA(wr_data_i[31:16]),
    .WE(wr_en_i),
    .MASK(16'h0000) );

SB_RAM40_4K #(
    .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .WRITE_MODE(0),
    .READ_MODE(0)
) ram256x16_q_inst (
    .RDATA(rd_data_o[15:0]),
    .RADDR(rd_addr),
    .RCLK(rd_clk_i),
    .RCLKE(1),    //<<
    .RE(rd_en_i),
    .WADDR(wr_addr),
    .WCLK (wr_clk_i),
    .WCLKE(wr_en_i),    //<<
    .WDATA(wr_data_i[15:0]),
    .WE(wr_en_i),
    .MASK(16'h0000) );

endmodule*/
